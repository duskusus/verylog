typedef logic[15:0] vec2[2];
typedef logic[15:0] vec3[3];
typedef logic[15:0] vec4[4];