`timescale 1ns / 1ps

module rasterizer(

    input logic Clk,
    
    // to framebuffer

    // from vertex memory

    
);

endmodule
