`timescale 1ns / 1ps

module rasterizer_control_unit(
    input logic Clk,
    
);

endmodule